.title KiCad schematic
JP1 /LV4 /LV3 GND 3.3V /LV2 /LV1 M06SIP
JP2 /A8 /A9 5V GND /HV3 /HV4 M06SIP
J5 3.3V GND /LV4 /LV3 NC_01 NC_02 3.3V NC_03 gyro connector
J3/J1 3.3V NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 5V GND NC_13 NC_14 /A9 /A8 NC_15 NC_16 NC_17 NC_18 ~
J2/J4 NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 NC_31 /HV4 /HV3 NC_32 NC_33 NC_34 NC_35 GND ~
U1 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 3.3V NC_42 NC_43 NC_44 NC_45 3.3V NC_46 NC_47 3.3V NC_48 GND /LV2 /LV1 NC_49 NC_50 NC_51 NC_52 NC_53 NC_54 NC_55 NC_56 NC_57 NC_58 NC_59 NodeMCU_1.0_(ESP-12E)
J1 /VIN GND /LV4 /LV3 /GPIO1 /XShutDown I2c
J4 7.5V GND Power supply
J2 /VIN GND /LV4 /LV3 /GPIO1 /XShutDown I2c
J3 /VIN GND /LV4 /LV3 /GPIO1 /XShutDown I2c
.end
